//ROM file for : bar_animation/bar_animation.hack
module hack_rom32k(clock, addr, out);
	input wire clock;
	input wire [14:0] addr;
	output reg [15:0] out;
	always @(posedge clock)
	begin
		case(addr)
			15'd00000 : out <= 16'b0000000000000000;
			15'd00001 : out <= 16'b1110110000010000;
			15'd00002 : out <= 16'b0000000000010000;
			15'd00003 : out <= 16'b1110001100001000;
			15'd00004 : out <= 16'b0001111101000000;
			15'd00005 : out <= 16'b1110110000010000;
			15'd00006 : out <= 16'b0000000000010001;
			15'd00007 : out <= 16'b1110001100001000;
			15'd00008 : out <= 16'b0100000000000000;
			15'd00009 : out <= 16'b1110110000010000;
			15'd00010 : out <= 16'b0000000000010000;
			15'd00011 : out <= 16'b1111000010010000;
			15'd00012 : out <= 16'b1110001100100000;
			15'd00013 : out <= 16'b1110101010001000;
			15'd00014 : out <= 16'b0000000000100001;
			15'd00015 : out <= 16'b1110110000010000;
			15'd00016 : out <= 16'b0000000000010000;
			15'd00017 : out <= 16'b1111000010001000;
			15'd00018 : out <= 16'b0100000000000000;
			15'd00019 : out <= 16'b1110110000010000;
			15'd00020 : out <= 16'b0000000000010000;
			15'd00021 : out <= 16'b1111000010010000;
			15'd00022 : out <= 16'b1110001100100000;
			15'd00023 : out <= 16'b1110111010001000;
			15'd00024 : out <= 16'b0000000000011110;
			15'd00025 : out <= 16'b1110110000010000;
			15'd00026 : out <= 16'b0000000000010010;
			15'd00027 : out <= 16'b1110001100001000;
			15'd00028 : out <= 16'b0000000000101010;
			15'd00029 : out <= 16'b1110101010000111;
			15'd00030 : out <= 16'b0000000000010001;
			15'd00031 : out <= 16'b1111110000010000;
			15'd00032 : out <= 16'b0000000000010000;
			15'd00033 : out <= 16'b1111010011010000;
			15'd00034 : out <= 16'b0000000000100110;
			15'd00035 : out <= 16'b1110001100000011;
			15'd00036 : out <= 16'b0000000000010000;
			15'd00037 : out <= 16'b1110101010001000;
			15'd00038 : out <= 16'b0000000000010001;
			15'd00039 : out <= 16'b1111110010001000;
			15'd00040 : out <= 16'b0000000000001000;
			15'd00041 : out <= 16'b1110101010000111;
			15'd00042 : out <= 16'b0111111111111111;
			15'd00043 : out <= 16'b1110110000010000;
			15'd00044 : out <= 16'b0000000000000000;
			15'd00045 : out <= 16'b1110001100001000;
			15'd00046 : out <= 16'b1110101010010000;
			15'd00047 : out <= 16'b0000000000110011;
			15'd00048 : out <= 16'b1110011111010010;
			15'd00049 : out <= 16'b0000000000101111;
			15'd00050 : out <= 16'b1110101010000111;
			15'd00051 : out <= 16'b0111111111111111;
			15'd00052 : out <= 16'b1110110000010000;
			15'd00053 : out <= 16'b0000000000000000;
			15'd00054 : out <= 16'b1111000010011000;
			15'd00055 : out <= 16'b0000000000010010;
			15'd00056 : out <= 16'b1111110000100000;
			15'd00057 : out <= 16'b1110001100000011;
			15'd00058 : out <= 16'b0000000000101110;
			15'd00059 : out <= 16'b1110101010000111;
			default:out <= 16'h0000;
		endcase
	end
endmodule
