
module hack_rom32k(clock, addr, out);

    input  wire         clock;
    input  wire [14:0]  addr;

    output reg  [15:0] out;

    always @(posedge clock)
    begin
        case(addr)
            // 15'h0000:out <= 16'b0101010101010101;
            // 15'h0001:out <= 16'b1110110000010000;
            // 15'h0002:out <= 16'b0100000000000000;
            // 15'h0003:out <= 16'b1110001100001000;
            // 15'h0004:out <= 16'b0000000000000100;
            // 15'h0005:out <= 16'b1110101010000111;
            // 15'h0006:out <= 16'b0000000000101000;
            // 15'h0007:out <= 16'b1110001100001000;
            // 15'h0008:out <= 16'b0000000000001000;
            // 15'h0009:out <= 16'b1110101010000111;
            // 15'h000a:out <= 16'b0000000000000000;
            // 15'h000b:out <= 16'b0000000000000000;
            15'd0000:out <= 16'b0000000001010101;
            15'd0001:out <= 16'b1110110000010000;
            15'd0002:out <= 16'b0100000000000000;
            15'd0003:out <= 16'b1110001100001000;
            15'd0004:out <= 16'b0000000000001010;
            15'd0005:out <= 16'b1110110000010000;
            15'd0006:out <= 16'b0000000000000001;
            15'd0007:out <= 16'b1110001100001000;
            15'd0008:out <= 16'b0000000000010100;
            15'd0009:out <= 16'b1110101010000111;
            15'd0010:out <= 16'b0000000010101010;
            15'd0011:out <= 16'b1110110000010000;
            15'd0012:out <= 16'b0100000000000000;
            15'd0013:out <= 16'b1110001100001000;
            15'd0014:out <= 16'b0000000000000000;
            15'd0015:out <= 16'b1110110000010000;
            15'd0016:out <= 16'b0000000000000001;
            15'd0017:out <= 16'b1110001100001000;
            15'd0018:out <= 16'b0000000000010100;
            15'd0019:out <= 16'b1110101010000111;
            15'd0020:out <= 16'b0111111111111111;
            15'd0021:out <= 16'b1110110000010000;
            15'd0022:out <= 16'b0000000000000000;
            15'd0023:out <= 16'b1110001100001000;
            15'd0024:out <= 16'b1110101010010000;
            15'd0025:out <= 16'b0000000000011101;
            15'd0026:out <= 16'b1110011111010010;
            15'd0027:out <= 16'b0000000000011001;
            15'd0028:out <= 16'b1110101010000111;
            15'd0029:out <= 16'b0010011100010000;
            15'd0030:out <= 16'b1110110000010000;
            15'd0031:out <= 16'b0000000000000000;
            15'd0032:out <= 16'b1111000010011000;
            15'd0033:out <= 16'b0000000000000001;
            15'd0034:out <= 16'b1111110000100000;
            15'd0035:out <= 16'b1110001100000011;
            15'd0036:out <= 16'b0000000000011000;
            15'd0037:out <= 16'b1110101010000111;
            default:out  <= 16'h0000;
        endcase
    end
endmodule
